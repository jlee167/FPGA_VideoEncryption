/*
Author: Jihoon Lee, Zachary Splingaire
Date: 5/8/2016
Module: quadMap
Function :	80 bit Key encryption through QuadMap Algorithm

Input: 80 bit key
output : Encryptiod 80 bit key
*/

module quadMap(input 						Clk,
													Reset,
													Run,
					 input [79:0]				in,
					 output logic [79:0]		out,
					 output						done);
		
endmodule 