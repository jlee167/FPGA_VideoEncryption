/*
IGNORE THIS FILE
Used for saving changed codes we are not sure about completely discarding 
*/