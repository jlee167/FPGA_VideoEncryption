/*
Author: Jihoon Lee, Zachary Splingaire
Date: 5/8/2016
Module: Unused Test Bench
*/



module testbench_test2();
/*
timeunit 10ns;

timeprecision 1ns;

logic Clk, Reset,	Cam_vsync, Cam_href, Cam_pclk;
logic [7:0]	Cam_data;
logic Cam_xclk, Cam_pwdn, Cam_reset_N, Cam_sdioc;
logic Cam_sdiod;

logic [7:0]  VGA_R, VGA_G, VGA_B;
logic VGA_CLK, VGA_SYNC_N, VGA_BLANK_N, VGA_VS, VGA_HS;

test2 test(.*);

always begin: CLOCK
	#1 Clk = ~Clk;
end

always begin: CAM_VSYNC
	#9408 Cam_vsync = 0;
	#1589952 Cam_vsync = 1;
end

always begin: CAM_href
	#62720 Cam_href = 1'b1;
	
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;
	#576 Cam_href = 1'b1;
	#2560 Cam_href = 1'b0;

	#31360 Cam_href = 1'b0;
	
end 

always begin: PIXEL_CLK
	#2 Cam_pclk = ~Cam_pclk;
end 

always begin: CAM_data
	#4 Cam_data = 8'b00010101;
	#4 Cam_data = 8'b01111100;
end 

initial begin
	Clk = 0;
	Cam_vsync = 1;
	Cam_href = 0;
	Cam_pclk = 0;
end

initial begin
	Reset = 1'b1;
	
	#2 Reset = 1'b0;
	
	#2 Reset = 1'b1;

	#15899520 Reset = 1'b0;
end */
endmodule 