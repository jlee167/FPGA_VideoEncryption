/*
Author: Jihoon Lee
Date: 3/8/2018
Module: LogicticMap
Function :	80 bit Key encryption through Logistic Map Algorithm

Input: 80 bit key
output : Encryptiod 80 bit key
*/

module logisticMap(input 						Clk,
														Reset,
														Run,
						 input [79:0]				in,
						 output logic [79:0]		out,
						 output						done);
			

			
endmodule 