/*
Author: Jihoon Lee, Zachary Splingaire
Date: 5/8/2016
Module: Multiplier80
Function :	Simple 80 bit Multiplication module
Input: 80 bit key
output : Encryptiod 80 bit key
*/

module multiplier80(input 						Clk,
														Reset,
														Run,
						  input [79:0] 			num1,
														num2,
						  output						done,
						  output logic [79:0]	out);
			
			
endmodule 